library verilog;
use verilog.vl_types.all;
entity test_vedic_8 is
end test_vedic_8;
